/mnt/c/users/dhava/Desktop/Web-dev/analog-clock